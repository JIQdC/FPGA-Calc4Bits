--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:08:47 08/15/2018
-- Design Name:   
-- Module Name:   C:/Documents and Settings/Solchu/My Documents/Projects/Calc4Bits/multtest.vhd
-- Project Name:  Calc4Bits
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: mult_sig_mag
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values\

USE ieee.numeric_std.ALL;
 
ENTITY multtest IS
END multtest;
 
ARCHITECTURE behavior OF multtest IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT mult_sig_mag
    PORT(
         a : IN  std_logic_vector(3 downto 0);
         b : IN  std_logic_vector(3 downto 0);
         mult : OUT  std_logic_vector(4 downto 0);
         over : OUT  std_logic
        );
    END COMPONENT;
    

   --Inputs
   signal a : std_logic_vector(3 downto 0) := (others => '0');
   signal b : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal mult : std_logic_vector(4 downto 0);
   signal over : std_logic;
	signal asig, bsig : std_logic;

 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: mult_sig_mag PORT MAP (
          a => a,
          b => b,
          mult => mult,
          over => over
        );
 

   -- Stimulus process
   stim_proc: process
   begin		
	--hago un doble loop de valores de a y b
	for avar in -7 to 7 loop
		--convierto el valor de avar en sig-mag y guardo el signo en asig
		if avar < 0 then
			a <= '1'& std_logic_vector(to_unsigned(abs(avar),3));
			asig <= '1';
		else 
			a <= '0'& std_logic_vector(to_unsigned(avar,3));
			asig <= '0';
		end if;
		
		for bvar in -7 to 7 loop
			--convierto el valor de bvar en sig-mag
			if bvar < 0 then
				b <= '1'& std_logic_vector(to_unsigned(abs(bvar),3));
				bsig <= '1';
			else 
				b <= '0'& std_logic_vector(to_unsigned(bvar,3));
				bsig <= '0';
			end if;
		
			--espero que ocurra la magia (?)
			wait for 1 ns;
			
			--primero chequeo que no haya hecho overflow (en cuyo caso no chequeo nada mas)
			if abs(avar*bvar) > 15 then
				assert over = '1' report "no hizo overflow" severity failure;
			--luego chequeo que no haga overflow, que la magnitud de la multiplicacion este bien y que el signo sea correcto
			else
				assert over = '0' report "hizo overflow cuando no deberia" severity failure;
				assert mult(3 downto 0)=std_logic_vector(to_unsigned(abs(avar*bvar),4)) report "magnitud de la mult esta mal" severity failure;
				assert mult(4)=(asig xor bsig) report "signo de la mult esta mal";
			end if;

		end loop;
	
	end loop;
	
	--aca respiramos nuevamente
	assert false report "todo bien :D" severity failure;
 
 
   end process;

END;
